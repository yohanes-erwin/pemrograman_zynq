`timescale 1ns / 1ps

module systolic_tb();
    localparam T = 10;
    
    reg clk;
    reg rst_n;
    reg en;
    reg clr;
    reg signed [15:0] a0, a1, a2, a3, a4, a5;
    reg in_valid;
    reg signed [15:0] b00, b01, b02, b03, b04, b05;
    reg signed [15:0] b10, b11, b12, b13, b14, b15;
    reg signed [15:0] b20, b21, b22, b23, b24, b25;
    reg signed [15:0] b30, b31, b32, b33, b34, b35;
    reg signed [15:0] b40, b41, b42, b43, b44, b45;
    reg signed [15:0] b50, b51, b52, b53, b54, b55;
    wire signed [15:0] y0, y1, y2, y3, y4, y5;
    wire out_valid;

    systolic
    #(
        .WIDTH(16),
        .FRAC_BIT(10)
    )
    dut
    (
        .clk(clk),
        .rst_n(rst_n),
        .en(en),
        .clr(clr),
        .a0(a0), .a1(a1), .a2(a2), .a3(a3), .a4(a4), .a5(a5),
        .in_valid(in_valid),
        .b00(b00), .b01(b01), .b02(b02), .b03(b03), .b04(b04), .b05(b05),
        .b10(b10), .b11(b11), .b12(b12), .b13(b13), .b14(b14), .b15(b15),
        .b20(b20), .b21(b21), .b22(b22), .b23(b23), .b24(b24), .b25(b25),
        .b30(b30), .b31(b31), .b32(b32), .b33(b33), .b34(b34), .b35(b35),
        .b40(b40), .b41(b41), .b42(b42), .b43(b43), .b44(b44), .b45(b45),
        .b50(b50), .b51(b51), .b52(b52), .b53(b53), .b54(b54), .b55(b55),
        .y0(y0), .y1(y1), .y2(y2), .y3(y3), .y4(y4), .y5(y5),
        .out_valid(out_valid)
    );

    always
    begin
        clk = 0;
        #(T/2);
        clk = 1;
        #(T/2);
    end

    initial
    begin
        en = 1;
        clr = 0;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0;
        in_valid = 0;
        b00 = 0; b01 = 0; b02 = 0; b03 = 0;  b04 = 0; b05 = 0;
        b10 = 0; b11 = 0; b12 = 0; b13 = 0;  b14 = 0; b15 = 0;
        b20 = 0; b21 = 0; b22 = 0; b23 = 0;  b24 = 0; b25 = 0;
        b30 = 0; b31 = 0; b32 = 0; b33 = 0;  b34 = 0; b35 = 0;
        b40 = 0; b41 = 0; b42 = 0; b43 = 0;  b44 = 0; b45 = 0;
        b50 = 0; b51 = 0; b52 = 0; b53 = 0;  b54 = 0; b55 = 0;
        
        rst_n = 0;
        #(T*5);
        rst_n = 1;
        #(T*5);
        
        // *** Testvector hidden layer 1 ***
        /*
         a = -1.2  1.3  1.7 -1.3 -1.3
              0.3  0.5  0.2  1   -1
              0.6  0.1  0.8  1.5 -1
              1.3 -1.2 -1.4  1.3 -0.9
              1.3  0.3  0.5  0.4 -1
        */
        /*
         b = 2  7 6 3  6 3
             10 2 8 10 9 2
             5  3 1 3  5 6
             3  3 6 1  6 10
             1  1 1 1  1 1
        */
        /*
         a*b =   13.9 -5.9  -4.2  11.9  3.9 -5.1
                 8.6   5.7  11     6.5 12.3 12.1
                 9.7  10.3  13.2   5.7 16.5 20.8
               -13.4   5.5   3.7 -11.9 -3.1  5.2
                8.3   11.4  12.1   7.8 14.4 10.5
        */
        b00 = 16'b000010_0000000000;  b01 = 16'b000111_0000000000;  b02 = 16'b000110_0000000000;  b03 = 16'b000011_0000000000; b04 = 16'b000110_0000000000; b05 = 16'b000011_0000000000;
        b10 = 16'b001010_0000000000;  b11 = 16'b000010_0000000000;  b12 = 16'b001000_0000000000;  b13 = 16'b001010_0000000000; b14 = 16'b001001_0000000000; b15 = 16'b000010_0000000000;
        b20 = 16'b000101_0000000000;  b21 = 16'b000011_0000000000;  b22 = 16'b000001_0000000000;  b23 = 16'b000011_0000000000; b24 = 16'b000101_0000000000; b25 = 16'b000110_0000000000;
        b30 = 16'b000011_0000000000;  b31 = 16'b000011_0000000000;  b32 = 16'b000110_0000000000;  b33 = 16'b000001_0000000000; b34 = 16'b000110_0000000000; b35 = 16'b001010_0000000000;
        b40 = 16'b000001_0000000000;  b41 = 16'b000001_0000000000;  b42 = 16'b000001_0000000000;  b43 = 16'b000001_0000000000; b44 = 16'b000001_0000000000; b45 = 16'b000001_0000000000;
        in_valid = 1;
        a0 = 16'b1111101100110011; a1 = 16'b0000010100110011; a2 = 16'b0000011011001100; a3 = 16'b1111101011001100; a4 = 16'b1111101011001100; a5 = 0;
        #T;
        a0 = 16'b0000000100110011; a1 = 16'b0000001000000000; a2 = 16'b0000000011001100; a3 = 16'b0000010000000000; a4 = 16'b1111110000000000; a5 = 0;
        #T;
        a0 = 16'b0000001001100110; a1 = 16'b0000000001100110; a2 = 16'b0000001100110011; a3 = 16'b0000011000000000; a4 = 16'b1111110000000000; a5 = 0;
        #T;
        a0 = 16'b0000010100110011; a1 = 16'b1111101100110011; a2 = 16'b1111101001100110; a3 = 16'b0000010100110011; a4 = 16'b1111110001100110; a5 = 0;
        #T;
        a0 = 16'b0000010100110011; a1 = 16'b0000000100110011; a2 = 16'b0000001000000000; a3 = 16'b0000000110011001; a4 = 16'b1111110000000000; a5 = 0;
        #T;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0;
        #T;
        in_valid = 0;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0;
        #(T*11);
        b00 = 0; b01 = 0; b02 = 0; b03 = 0;  b04 = 0; b05 = 0;
        b10 = 0; b11 = 0; b12 = 0; b13 = 0;  b14 = 0; b15 = 0;
        b20 = 0; b21 = 0; b22 = 0; b23 = 0;  b24 = 0; b25 = 0;
        b30 = 0; b31 = 0; b32 = 0; b33 = 0;  b34 = 0; b35 = 0;
        b40 = 0; b41 = 0; b42 = 0; b43 = 0;  b44 = 0; b45 = 0;
        b50 = 0; b51 = 0; b52 = 0; b53 = 0;  b54 = 0; b55 = 0;
        #(T*10);
        
        // *** Testvector hidden layer 2 ***
        /*
         a =  5.2 -0.3 0.8 -3.5 0.1	-1.5
             -4.8  0.1 0.7  4	0.9	-1.4
        */
        /*
         b = 1 0 0 1 1 0
             1 1 1 1 1 1
             1 1 1 1 1 1
             0 1 1 0 0 1
             1 1 1 1 1 1
             1 1 1 1 1 1
        */
        /*
         a*b =  4.29 -4.37 -4.23 4.29 4.04 -4.34
               -4.50 4.27 4.13 -4.50 -4.23 4.24
        */
        b00 = 16'b000001_0000000000;  b01 = 16'b000000_0000000000;  b02 = 16'b000000_0000000000;  b03 = 16'b000001_0000000000; b04 = 16'b000001_0000000000; b05 = 16'b000000_0000000000;
        b10 = 16'b000001_0000000000;  b11 = 16'b000001_0000000000;  b12 = 16'b000001_0000000000;  b13 = 16'b000001_0000000000; b14 = 16'b000001_0000000000; b15 = 16'b000001_0000000000;
        b20 = 16'b000001_0000000000;  b21 = 16'b000001_0000000000;  b22 = 16'b000001_0000000000;  b23 = 16'b000001_0000000000; b24 = 16'b000001_0000000000; b25 = 16'b000001_0000000000;
        b30 = 16'b000000_0000000000;  b31 = 16'b000001_0000000000;  b32 = 16'b000001_0000000000;  b33 = 16'b000000_0000000000; b34 = 16'b000000_0000000000; b35 = 16'b000001_0000000000;
        b40 = 16'b000001_0000000000;  b41 = 16'b000001_0000000000;  b42 = 16'b000001_0000000000;  b43 = 16'b000001_0000000000; b44 = 16'b000001_0000000000; b45 = 16'b000001_0000000000;
        b50 = 16'b000001_0000000000;  b51 = 16'b000001_0000000000;  b52 = 16'b000001_0000000000;  b53 = 16'b000001_0000000000; b54 = 16'b000001_0000000000; b55 = 16'b000001_0000000000;
        in_valid = 1;
        a0 = 16'b0001010011001100; a1 = 16'b1111111011001100; a2 = 16'b0000001100110011; a3 = 16'b1111001000000000; a4 = 16'b0000000001100110; a5 = 16'b1111101000000000;
        #T;
        a0 = 16'b1110110011001100; a1 = 16'b0000000001100110; a2 = 16'b0000001011001100; a3 = 16'b0001000000000000; a4 = 16'b0000001110011001; a5 = 16'b1111101001100110;
        #T;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0;
        #T;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0;
        #T;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0;
        #T;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0;
        #T;
        in_valid = 0;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0;
        #(T*11);
        b00 = 0; b01 = 0; b02 = 0; b03 = 0;  b04 = 0; b05 = 0;
        b10 = 0; b11 = 0; b12 = 0; b13 = 0;  b14 = 0; b15 = 0;
        b20 = 0; b21 = 0; b22 = 0; b23 = 0;  b24 = 0; b25 = 0;
        b30 = 0; b31 = 0; b32 = 0; b33 = 0;  b34 = 0; b35 = 0;
        b40 = 0; b41 = 0; b42 = 0; b43 = 0;  b44 = 0; b45 = 0;
        b50 = 0; b51 = 0; b52 = 0; b53 = 0;  b54 = 0; b55 = 0;
        #(T*10);
    end

endmodule
