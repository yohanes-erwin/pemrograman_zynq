// *** Author : Erwin Ouyang
// *** Date   : 10 May 2018
`timescale 1ns / 1ps

module matrix_dp_tb();
    localparam T = 10;
    
    reg clk;
    reg rst_n;
    reg en;
    reg clr;
    reg signed [15:0] x0, x1, x2, x3, x4, x5, x6, x7;
    reg signed [15:0] w00, w01, w02, w03, w04, w05, w06, w07;
    reg signed [15:0] w10, w11, w12, w13, w14, w15, w16, w17;
    reg signed [15:0] w20, w21, w22, w23, w24, w25, w26, w27;
    reg signed [15:0] w30, w31, w32, w33, w34, w35, w36, w37;
    reg signed [15:0] w40, w41, w42, w43, w44, w45, w46, w47;
    reg signed [15:0] w50, w51, w52, w53, w54, w55, w56, w57;
    reg signed [15:0] w60, w61, w62, w63, w64, w65, w66, w67;
    reg signed [15:0] w70, w71, w72, w73, w74, w75, w76, w77;
    wire signed [15:0] z0, z1, z2, z3, z4, z5, z6, z7;

    matrix_dp uut
    (
        .clk(clk),
        .rst_n(rst_n),
        .en(en),
        .clr(clr),
        .x0(x0), .x1(x1), .x2(x2), .x3(x3), .x4(x4), .x5(x5), .x6(x6), .x7(x7),
        .w00(w00), .w01(w01), .w02(w02), .w03(w03), .w04(w04), .w05(w05), .w06(w06), .w07(w07),
        .w10(w10), .w11(w11), .w12(w12), .w13(w13), .w14(w14), .w15(w15), .w16(w16), .w17(w17),
        .w20(w20), .w21(w21), .w22(w22), .w23(w23), .w24(w24), .w25(w25), .w26(w26), .w27(w27),
        .w30(w30), .w31(w31), .w32(w32), .w33(w33), .w34(w34), .w35(w35), .w36(w36), .w37(w37),
        .w40(w40), .w41(w41), .w42(w42), .w43(w43), .w44(w44), .w45(w45), .w46(w46), .w47(w47),
        .w50(w50), .w51(w51), .w52(w52), .w53(w53), .w54(w54), .w55(w55), .w56(w56), .w57(w57),
        .w60(w60), .w61(w61), .w62(w62), .w63(w63), .w64(w64), .w65(w65), .w66(w66), .w67(w67),
        .w70(w70), .w71(w71), .w72(w72), .w73(w73), .w74(w74), .w75(w75), .w76(w76), .w77(w77),
        .z0(z0), .z1(z1), .z2(z2), .z3(z3), .z4(z4), .z5(z5), .z6(z6), .z7(z7)
    );

    always
    begin
        clk = 0;
        #(T/2);
        clk = 1;
        #(T/2);
    end

    initial
    begin
        rst_n = 0;
        en = 0;
        clr = 0;
        x0 = 0; x1 = 0; x2 = 0; x3 = 0; x4 = 0; x5 = 0; x6 = 0; x7 = 0;
        w00 = 0; w01 = 0; w02 = 0; w03 = 0; w04 = 0; w05 = 0; w06 = 0; w07 = 0;
        w10 = 0; w11 = 0; w12 = 0; w13 = 0; w14 = 0; w15 = 0; w16 = 0; w17 = 0;
        w20 = 0; w21 = 0; w22 = 0; w23 = 0; w24 = 0; w25 = 0; w26 = 0; w27 = 0;
        w30 = 0; w31 = 0; w32 = 0; w33 = 0; w34 = 0; w35 = 0; w36 = 0; w37 = 0;
        w40 = 0; w41 = 0; w42 = 0; w43 = 0; w44 = 0; w45 = 0; w46 = 0; w47 = 0;
        w50 = 0; w51 = 0; w52 = 0; w53 = 0; w54 = 0; w55 = 0; w56 = 0; w57 = 0;
        w60 = 0; w61 = 0; w62 = 0; w63 = 0; w64 = 0; w65 = 0; w66 = 0; w67 = 0;
        w70 = 0; w71 = 0; w72 = 0; w73 = 0; w74 = 0; w75 = 0; w76 = 0; w77 = 0;
        #(T*5);
        rst_n = 1;
        en = 1;
        #(T*5);
        
        w00 = 16'b00_0010_0001_1001_10; w01 = 16'b00_0001_1000_0110_01; w02 = 16'b00_0000_1110_0000_00;
        w10 = 16'b00_0000_1000_0111_00; w11 = 16'b00_0010_1100_0000_01; w12 = 16'b00_0001_1000_1100_00;
        w20 = 16'b00_0011_1110_010_00; w21 = 16'b00_0100_110_0001_00; w22 = 16'b00_0000_1000_0100_11;
        
        x0 = 16'b00_0001_1000_0010_10; x1 = 0; x2 = 0;
        #T;
        x0 = 16'b00_0011_1110_0110_10; x1 = 16'b00_0010_1010_0000_00; x2 = 0;
        #T;
        x0 = 16'b00_0000_1111_0000_11; x1 = 16'b00_0001_1000_0000_11; x2 = 16'b00_0000_1111_1111_00;
        #T;
        x0 = 0; x1 = 16'b00_0000_1010_0000_00; x2 = 16'b00_0000_1000_0000_00;
        #T;
        x0 = 0; x1 = 0; x2 = 16'b00_0000_1000_0101_00;
        #T;
        x0 = 0; x1 = 0; x2 = 0;
        #T;
    end

endmodule
