`timescale 1ns / 1ps

module systolic_nn_tb();
    localparam T = 10;
    
    reg clk;
    reg rst_n;
    reg en;
    reg clr;
    reg signed [15:0] a0, a1, a2, a3;
    reg in_valid;
    reg signed [15:0] b00, b01, b02, b03;
    reg signed [15:0] b10, b11, b12, b13;
    reg signed [15:0] b20, b21, b22, b23;
    reg signed [15:0] b30, b31, b32, b33;
    wire signed [15:0] y0, y1, y2, y3;
    wire out_valid;

    systolic
    #(
        .WIDTH(16),
        .FRAC_BIT(10)
    )
    dut
    (
        .clk(clk),
        .rst_n(rst_n),
        .en(en),
        .clr(clr),
        .a0(a0), .a1(a1), .a2(a2), .a3(a3),
        .in_valid(in_valid),
        .b00(b00), .b01(b01), .b02(b02), .b03(b03),
        .b10(b10), .b11(b11), .b12(b12), .b13(b13),
        .b20(b20), .b21(b21), .b22(b22), .b23(b23),
        .b30(b30), .b31(b31), .b32(b32), .b33(b33),
        .y0(y0), .y1(y1), .y2(y2), .y3(y3),
        .out_valid(out_valid)
    );

    always
    begin
        clk = 0;
        #(T/2);
        clk = 1;
        #(T/2);
    end

    initial
    begin
        en = 1;
        clr = 0;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0;
        in_valid = 0;
        b00 = 0; b01 = 0; b02 = 0; b03 = 0;
        b10 = 0; b11 = 0; b12 = 0; b13 = 0;
        b20 = 0; b21 = 0; b22 = 0; b23 = 0;
        b30 = 0; b31 = 0; b32 = 0; b33 = 0;
        
        rst_n = 0;
        #(T*5);
        rst_n = 1;
        #(T*5);
 
        // *** Testvector 1 ***
        /*
         a = 1.37    1.37  -19.88
             0.77    0.97   -0.90
             1.05    0.64   -0.89
        */
        /*
         b = 8     8     5     5
             8     5     8     5
             1     1     1     1
        */
        /*
         a*b =  2.04   -2.07   -2.07   -6.18
               13.02   10.11   10.71    7.80
               12.63   10.71    9.48    7.56
        */
        b00 = 16'b0010000000000000;  b01 = 16'b0010000000000000;  b02 = 16'b0001010000000000;  b03 = 16'b0001010000000000;
        b10 = 16'b0010000000000000;  b11 = 16'b0001010000000000;  b12 = 16'b0010000000000000;  b13 = 16'b0001010000000000;
        b20 = 16'b0000010000000000;  b21 = 16'b0000010000000000;  b22 = 16'b0000010000000000;  b23 = 16'b0000010000000000;
        b30 = 0;  b31 = 0;  b32 = 0;  b33 = 0;
        in_valid = 1;
        a0 = 16'b0000010101111010; a1 = 16'b0000010101111010; a2 = 16'b1011000001111010; a3 = 0;
        #T;
        a0 = 16'b0000001100010100; a1 = 16'b0000001111100001; a2 = 16'b1111110001100110; a3 = 0;
        #T;
        a0 = 16'b0000010000110011; a1 = 16'b0000001010001111; a2 = 16'b1111110001110000; a3 = 0;
        #T;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0;
        #T;
        in_valid = 0;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0;
        #(T*7);
        b00 = 0; b01 = 0; b02 = 0; b03 = 0;
        b10 = 0; b11 = 0; b12 = 0; b13 = 0;
        b20 = 0; b21 = 0; b22 = 0; b23 = 0;
        b30 = 0; b31 = 0; b32 = 0; b33 = 0;
 
        // *** Testvector 2 ***
        /*
         a =  7.11   -1.31    0.08   -2.59
             -7.10    1.63    1.97    0.20
        */
        /*
         b = 0.8849    0.1120    0.1120    0.0021
             1.0000    1.0000    1.0000    0.9996
             1.0000    1.0000    0.9999    0.9995
             1.0000    1.0000    1.0000    1.0000
        */
        /*
         a*b =  2.4719   -3.0233   -3.0233   -3.8048
               -2.4830    3.0044    3.0043    3.7836
        */
        b00 = 16'b0000001110001010;  b01 = 16'b0000000001110010;  b02 = 16'b0000000001110010;  b03 = 16'b0000000000000010;
        b10 = 16'b0000010000000000;  b11 = 16'b0000010000000000;  b12 = 16'b0000010000000000;  b13 = 16'b0000001111111111;
        b20 = 16'b0000010000000000;  b21 = 16'b0000010000000000;  b22 = 16'b0000001111111111;  b23 = 16'b0000001111111111;
        b30 = 16'b0000010000000000;  b31 = 16'b0000010000000000;  b32 = 16'b0000010000000000;  b33 = 16'b0000010000000000;
        in_valid = 1;
        a0 = 16'b0001110001110000; a1 = 16'b1111101011000010; a2 = 16'b0000000001010001; a3 = 16'b1111010110100011;
        #T;
        a0 = 16'b1110001110011001; a1 = 16'b0000011010000101; a2 = 16'b0000011111100001; a3 = 16'b0000000011001100;
        #T;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0;
        #T;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0;
        #T;
        in_valid = 0;
        a0 = 0; a1 = 0; a2 = 0; a3 = 0;
        #(T*7);
        b00 = 0; b01 = 0; b02 = 0; b03 = 0;
        b10 = 0; b11 = 0; b12 = 0; b13 = 0;
        b20 = 0; b21 = 0; b22 = 0; b23 = 0;
        b30 = 0; b31 = 0; b32 = 0; b33 = 0;
    end

endmodule
